Library IEEE;
Use IEEE.Std_logic_1164.all;
--  Defines a design entity
package EvParity;
function Eparity (a:std_logic_vector(3 downto 0)) 

architecture behaviour of package is
begin
    process

    begin

        wait;
    end process;
end behaviour;
